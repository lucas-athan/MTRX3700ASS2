module grayscale_producer #(
    parameter WIDTH  = 640,
    parameter HEIGHT = 480
)(
    input  logic       clk,
    input  logic       reset,
    input  logic       ready,
    output logic [7:0] pixel_out,
    output logic       valid,
    output logic       startofpacket,
    output logic       endofpacket
);

    localparam int NUMPIXELS = WIDTH * HEIGHT;   // 307,200

    // Pixel counter
    logic [18:0] pixel_index;

    always_ff @(posedge clk) begin
        if (reset)
            pixel_index <= 19'd0;
        else if (valid && ready) begin
            if (pixel_index == NUMPIXELS-1)
                pixel_index <= 19'd0;
            else
                pixel_index <= pixel_index + 19'd1;
        end
    end

    // Instantiate ROM generated by MegaWizard
    wire [7:0] rom_q;

    ImageRom image_rom_inst (
        .address(pixel_index), // 19-bit address
        .clock(clk),           // same clock
        .q(rom_q)              // ROM output
    );

    // Outputs
    assign pixel_out     = rom_q;
    assign valid         = ~reset;
    assign startofpacket = (pixel_index == 0);
    assign endofpacket   = (pixel_index == NUMPIXELS-1);

endmodule
